
module incr_A(output [7:0] out, input [7:0] a);

assign out = a + 1;

endmodule